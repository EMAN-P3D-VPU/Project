////////////////////////////////////////////////////////////////////////////////
// execute.v
// Dan Wortmann
//
// Description:
// 
////////////////////////////////////////////////////////////////////////////////
module execute();
////////////
// Inputs /
//////////

/////////////
// Outputs /
///////////

/////////////////////////////
// Signals/Logic/Registers /
///////////////////////////

///////////////////
// Interconnects /
/////////////////

////////////////////////////////////////////////////////////////////////////////
// execute
////

// Memory R/W //

// Write Back Logic //

endmodule
