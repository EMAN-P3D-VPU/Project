
 
 
 




window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"


      waveform add -signals /frame_cell_block_tb/status
      waveform add -signals /frame_cell_block_tb/frame_cell_block_synth_inst/bmg_port/CLKA
      waveform add -signals /frame_cell_block_tb/frame_cell_block_synth_inst/bmg_port/ADDRA
      waveform add -signals /frame_cell_block_tb/frame_cell_block_synth_inst/bmg_port/DINA
      waveform add -signals /frame_cell_block_tb/frame_cell_block_synth_inst/bmg_port/WEA
      waveform add -signals /frame_cell_block_tb/frame_cell_block_synth_inst/bmg_port/DOUTA
console submit -using simulator -wait no "run"
