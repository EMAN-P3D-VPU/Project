//module checks the distances between testpoints and real point
//outputs which delt is closer to the real point
module delta_select(x_0, x_1, y_0, y_1, dy, );




endmodule
