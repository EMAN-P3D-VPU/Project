////////////////////////////////////////////////////////////////////////////////
// cpu_memory_control.v
// Dan Wortmann
//
// Description:
// 
////////////////////////////////////////////////////////////////////////////////
module cpu_memory_control();
////////////
// Inputs /
//////////

/////////////
// Outputs /
///////////

/////////////////////////////
// Signals/Logic/Registers /
///////////////////////////

///////////////////
// Interconnects /
/////////////////

////////////////////////////////////////////////////////////////////////////////
// cpu_memory_control
////

// Main CPU Memory //

// I-Cache //

// Cache Controller //

endmodule
