////////////////////////////////////////////////////////////////////////////////
// alu.v
// Dan Wortmann
//
// Description:
// 
////////////////////////////////////////////////////////////////////////////////
module alu();
////////////
// Inputs /
//////////

/////////////
// Outputs /
///////////

/////////////////////////////
// Signals/Logic/Registers /
///////////////////////////

///////////////////
// Interconnects /
/////////////////

////////////////////////////////////////////////////////////////////////////////
// alu
////

endmodule
