
module test(in, out);

input in;
output out;

reg x;

assign x = 2;

endmodule;