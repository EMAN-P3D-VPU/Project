////////////////////////////////////////////////////////////////////////////////
// cache.v
// Dan Wortmann
//
// Description:
// 
////////////////////////////////////////////////////////////////////////////////
module cache();
////////////
// Inputs /
//////////

/////////////
// Outputs /
///////////

/////////////////////////////
// Signals/Logic/Registers /
///////////////////////////

///////////////////
// Interconnects /
/////////////////

////////////////////////////////////////////////////////////////////////////////
// cache
////

endmodule
