module steep_calculator_TB ();

steep_calculator steep_calc(line_cap_reg, dy, dx, slope_steep);
endmodule