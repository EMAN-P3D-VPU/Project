////////////////////////////////////////////////////////////////////////////////
// memory_writeback.v
// Dan Wortmann
//
// Description:
// 
////////////////////////////////////////////////////////////////////////////////
module memory_writeback();
////////////
// Inputs /
//////////

/////////////
// Outputs /
///////////

/////////////////////////////
// Signals/Logic/Registers /
///////////////////////////

///////////////////
// Interconnects /
/////////////////

////////////////////////////////////////////////////////////////////////////////
// memory_writeback
////

// Memory R/W //

// Write Back Logic //

endmodule