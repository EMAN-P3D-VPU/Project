module frame_cell(
				// General Inputs
				input clk,

				// Writing
				input [9:0] write_frame_width,
				input [8:0] write_frame_height,
				input write_enable,
				input [2:0] write_data,

				// Reading
				input [9:0] read_frame_width,
				input [8:0] read_frame_height,
				output [2:0] read_data);

// simple dual port RAM with a common clock
// write width - 3
// write detph - 307200 (640 x 480)
// initialize everything to 0
frame_cell_block block_mem(
			.addra({write_frame_width, write_frame_height}),
			.dina(write_data),
			.wea(write_enable),
			.clka(clk),
			.addrb({read_frame_width, read_frame_height}),
			.clkb(clk),
			.doutb(read_data));

endmodule