////////////////////////////////////////////////////////////////////////////////
// instruction_decode_execute.v
// Dan Wortmann
//
// Description:
// 
////////////////////////////////////////////////////////////////////////////////
module instruction_decode_execute();
////////////
// Inputs /
//////////

/////////////
// Outputs /
///////////

/////////////////////////////
// Signals/Logic/Registers /
///////////////////////////

///////////////////
// Interconnects /
/////////////////

////////////////////////////////////////////////////////////////////////////////
// instruction_decode_execute
////

// Control //

// Register File //

// ALU //

// Branching Unit //

endmodule
