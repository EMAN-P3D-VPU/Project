////////////////////////////////////////////////////////////////////////////////
// instruction_decode.v
// Dan Wortmann
//
// Description:
// 
////////////////////////////////////////////////////////////////////////////////
module instruction_decode();
////////////
// Inputs /
//////////

/////////////
// Outputs /
///////////

/////////////////////////////
// Signals/Logic/Registers /
///////////////////////////

///////////////////
// Interconnects /
/////////////////

////////////////////////////////////////////////////////////////////////////////
// instruction_decode
////

// Control //

// Register File //

// ALU //

// Branching Unit //

endmodule
